`define TRACE_PORTAL 
`define ConnectalVersion 20.06.4
`define NumberOfMasters 1
`define PinType Empty
`define PinTypeInclude Misc
`define NumberOfUserTiles 1
`define SlaveDataBusWidth 32
`define SlaveControlAddrWidth 5
`define BurstLenSize 10
`define project_dir $(DTOP)
`define MainClockPeriod 20
`define DerivedClockPeriod 10.000000
`define CnocTop 
`define XsimHostInterface 
`define PhysAddrWidth 40
`define SIMULATION 
`define CONNECTAL_BITS_DEPENDENCES bsim
`define BOARD_bluesim 
